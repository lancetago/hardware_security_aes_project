-- Inverse Substitution Box VHDL module
-- LUT that stores the AES inverse S-Box
-- 

library ieee;
use ieee.std_logic_1164.all;

entity inv_s_box is
port (
    i_byte : in std_logic_vector(7 downto 0);
    o_byte : out std_logic_vector(7 downto 0)
);
end inv_s_box;

architecture behavioral of inv_s_box is

begin
	process (i_byte)
	begin
		case i_byte is
			when x"00" => o_byte <= x"52";
			when x"01" => o_byte <= x"09";
			when x"02" => o_byte <= x"6a";
			when x"03" => o_byte <= x"d5";
			when x"04" => o_byte <= x"30";
			when x"05" => o_byte <= x"36";
			when x"06" => o_byte <= x"a5";
			when x"07" => o_byte <= x"38";
			when x"08" => o_byte <= x"bf";
			when x"09" => o_byte <= x"40";
			when x"0a" => o_byte <= x"a3";
			when x"0b" => o_byte <= x"9e";
			when x"0c" => o_byte <= x"81";
			when x"0d" => o_byte <= x"f3";
			when x"0e" => o_byte <= x"d7";
			when x"0f" => o_byte <= x"fb";
			when x"10" => o_byte <= x"7c";
			when x"11" => o_byte <= x"e3";
			when x"12" => o_byte <= x"39";
			when x"13" => o_byte <= x"82";
			when x"14" => o_byte <= x"9b";
			when x"15" => o_byte <= x"2f";
			when x"16" => o_byte <= x"ff";
			when x"17" => o_byte <= x"87";
			when x"18" => o_byte <= x"34";
			when x"19" => o_byte <= x"8e";
			when x"1a" => o_byte <= x"43";
			when x"1b" => o_byte <= x"44";
			when x"1c" => o_byte <= x"c4";
			when x"1d" => o_byte <= x"de";
			when x"1e" => o_byte <= x"e9";
			when x"1f" => o_byte <= x"cb";
			when x"20" => o_byte <= x"54";
			when x"21" => o_byte <= x"7b";
			when x"22" => o_byte <= x"94";
			when x"23" => o_byte <= x"32";
			when x"24" => o_byte <= x"a6";
			when x"25" => o_byte <= x"c2";
			when x"26" => o_byte <= x"23";
			when x"27" => o_byte <= x"3d";
			when x"28" => o_byte <= x"ee";
			when x"29" => o_byte <= x"4c";
			when x"2a" => o_byte <= x"95";
			when x"2b" => o_byte <= x"0b";
			when x"2c" => o_byte <= x"42";
			when x"2d" => o_byte <= x"fa";
			when x"2e" => o_byte <= x"c3";
			when x"2f" => o_byte <= x"4e";
			when x"30" => o_byte <= x"08";
			when x"31" => o_byte <= x"2e";
			when x"32" => o_byte <= x"a1";
			when x"33" => o_byte <= x"66";
			when x"34" => o_byte <= x"28";
			when x"35" => o_byte <= x"d9";
			when x"36" => o_byte <= x"24";
			when x"37" => o_byte <= x"b2";
			when x"38" => o_byte <= x"76";
			when x"39" => o_byte <= x"5b";
			when x"3a" => o_byte <= x"a2";
			when x"3b" => o_byte <= x"49";
			when x"3c" => o_byte <= x"6d";
			when x"3d" => o_byte <= x"8b";
			when x"3e" => o_byte <= x"d1";
			when x"3f" => o_byte <= x"25";
			when x"40" => o_byte <= x"72";
			when x"41" => o_byte <= x"f8";
			when x"42" => o_byte <= x"f6";
			when x"43" => o_byte <= x"64";
			when x"44" => o_byte <= x"86";
			when x"45" => o_byte <= x"68";
			when x"46" => o_byte <= x"98";
			when x"47" => o_byte <= x"16";
			when x"48" => o_byte <= x"d4";
			when x"49" => o_byte <= x"a4";
			when x"4a" => o_byte <= x"5c";
			when x"4b" => o_byte <= x"cc";
			when x"4c" => o_byte <= x"5d";
			when x"4d" => o_byte <= x"65";
			when x"4e" => o_byte <= x"b6";
			when x"4f" => o_byte <= x"92";
			when x"50" => o_byte <= x"6c";
			when x"51" => o_byte <= x"70";
			when x"52" => o_byte <= x"48";
			when x"53" => o_byte <= x"50";
			when x"54" => o_byte <= x"fd";
			when x"55" => o_byte <= x"ed";
			when x"56" => o_byte <= x"b9";
			when x"57" => o_byte <= x"da";
			when x"58" => o_byte <= x"5e";
			when x"59" => o_byte <= x"15";
			when x"5a" => o_byte <= x"46";
			when x"5b" => o_byte <= x"57";
			when x"5c" => o_byte <= x"a7";
			when x"5d" => o_byte <= x"8d";
			when x"5e" => o_byte <= x"9d";
			when x"5f" => o_byte <= x"84";
			when x"60" => o_byte <= x"90";
			when x"61" => o_byte <= x"d8";
			when x"62" => o_byte <= x"ab";
			when x"63" => o_byte <= x"00";
			when x"64" => o_byte <= x"8c";
			when x"65" => o_byte <= x"bc";
			when x"66" => o_byte <= x"d3";
			when x"67" => o_byte <= x"0a";
			when x"68" => o_byte <= x"f7";
			when x"69" => o_byte <= x"e4";
			when x"6a" => o_byte <= x"58";
			when x"6b" => o_byte <= x"05";
			when x"6c" => o_byte <= x"b8";
			when x"6d" => o_byte <= x"b3";
			when x"6e" => o_byte <= x"45";
			when x"6f" => o_byte <= x"06";
			when x"70" => o_byte <= x"d0";
			when x"71" => o_byte <= x"2c";
			when x"72" => o_byte <= x"1e";
			when x"73" => o_byte <= x"8f";
			when x"74" => o_byte <= x"ca";
			when x"75" => o_byte <= x"3f";
			when x"76" => o_byte <= x"0f";
			when x"77" => o_byte <= x"02";
			when x"78" => o_byte <= x"c1";
			when x"79" => o_byte <= x"af";
			when x"7a" => o_byte <= x"bd";
			when x"7b" => o_byte <= x"03";
			when x"7c" => o_byte <= x"01";
			when x"7d" => o_byte <= x"13";
			when x"7e" => o_byte <= x"8a";
			when x"7f" => o_byte <= x"6b";
			when x"80" => o_byte <= x"3a";
			when x"81" => o_byte <= x"91";
			when x"82" => o_byte <= x"11";
			when x"83" => o_byte <= x"41";
			when x"84" => o_byte <= x"4f";
			when x"85" => o_byte <= x"67";
			when x"86" => o_byte <= x"dc";
			when x"87" => o_byte <= x"ea";
			when x"88" => o_byte <= x"97";
			when x"89" => o_byte <= x"f2";
			when x"8a" => o_byte <= x"cf";
			when x"8b" => o_byte <= x"ce";
			when x"8c" => o_byte <= x"f0";
			when x"8d" => o_byte <= x"b4";
			when x"8e" => o_byte <= x"e6";
			when x"8f" => o_byte <= x"73";
			when x"90" => o_byte <= x"96";
			when x"91" => o_byte <= x"ac";
			when x"92" => o_byte <= x"74";
			when x"93" => o_byte <= x"22";
			when x"94" => o_byte <= x"e7";
			when x"95" => o_byte <= x"ad";
			when x"96" => o_byte <= x"35";
			when x"97" => o_byte <= x"85";
			when x"98" => o_byte <= x"e2";
			when x"99" => o_byte <= x"f9";
			when x"9a" => o_byte <= x"37";
			when x"9b" => o_byte <= x"e8";
			when x"9c" => o_byte <= x"1c";
			when x"9d" => o_byte <= x"75";
			when x"9e" => o_byte <= x"df";
			when x"9f" => o_byte <= x"6e";
			when x"a0" => o_byte <= x"47";
			when x"a1" => o_byte <= x"f1";
			when x"a2" => o_byte <= x"1a";
			when x"a3" => o_byte <= x"71";
			when x"a4" => o_byte <= x"1d";
			when x"a5" => o_byte <= x"29";
			when x"a6" => o_byte <= x"c5";
			when x"a7" => o_byte <= x"89";
			when x"a8" => o_byte <= x"6f";
			when x"a9" => o_byte <= x"b7";
			when x"aa" => o_byte <= x"62";
			when x"ab" => o_byte <= x"0e";
			when x"ac" => o_byte <= x"aa";
			when x"ad" => o_byte <= x"18";
			when x"ae" => o_byte <= x"be";
			when x"af" => o_byte <= x"1b";
			when x"b0" => o_byte <= x"fc";
			when x"b1" => o_byte <= x"56";
			when x"b2" => o_byte <= x"3e";
			when x"b3" => o_byte <= x"4b";
			when x"b4" => o_byte <= x"c6";
			when x"b5" => o_byte <= x"d2";
			when x"b6" => o_byte <= x"79";
			when x"b7" => o_byte <= x"20";
			when x"b8" => o_byte <= x"9a";
			when x"b9" => o_byte <= x"db";
			when x"ba" => o_byte <= x"c0";
			when x"bb" => o_byte <= x"fe";
			when x"bc" => o_byte <= x"78";
			when x"bd" => o_byte <= x"cd";
			when x"be" => o_byte <= x"5a";
			when x"bf" => o_byte <= x"f4";
			when x"c0" => o_byte <= x"1f";
			when x"c1" => o_byte <= x"dd";
			when x"c2" => o_byte <= x"a8";
			when x"c3" => o_byte <= x"33";
			when x"c4" => o_byte <= x"88";
			when x"c5" => o_byte <= x"07";
			when x"c6" => o_byte <= x"c7";
			when x"c7" => o_byte <= x"31";
			when x"c8" => o_byte <= x"b1";
			when x"c9" => o_byte <= x"12";
			when x"ca" => o_byte <= x"10";
			when x"cb" => o_byte <= x"59";
			when x"cc" => o_byte <= x"27";
			when x"cd" => o_byte <= x"80";
			when x"ce" => o_byte <= x"ec";
			when x"cf" => o_byte <= x"5f";
			when x"d0" => o_byte <= x"60";
			when x"d1" => o_byte <= x"51";
			when x"d2" => o_byte <= x"7f";
			when x"d3" => o_byte <= x"a9";
			when x"d4" => o_byte <= x"19";
			when x"d5" => o_byte <= x"b5";
			when x"d6" => o_byte <= x"4a";
			when x"d7" => o_byte <= x"0d";
			when x"d8" => o_byte <= x"2d";
			when x"d9" => o_byte <= x"e5";
			when x"da" => o_byte <= x"7a";
			when x"db" => o_byte <= x"9f";
			when x"dc" => o_byte <= x"93";
			when x"dd" => o_byte <= x"c9";
			when x"de" => o_byte <= x"9c";
			when x"df" => o_byte <= x"ef";
			when x"e0" => o_byte <= x"a0";
			when x"e1" => o_byte <= x"e0";
			when x"e2" => o_byte <= x"3b";
			when x"e3" => o_byte <= x"4d";
			when x"e4" => o_byte <= x"ae";
			when x"e5" => o_byte <= x"2a";
			when x"e6" => o_byte <= x"f5";
			when x"e7" => o_byte <= x"b0";
			when x"e8" => o_byte <= x"c8";
			when x"e9" => o_byte <= x"eb";
			when x"ea" => o_byte <= x"bb";
			when x"eb" => o_byte <= x"3c";
			when x"ec" => o_byte <= x"83";
			when x"ed" => o_byte <= x"53";
			when x"ee" => o_byte <= x"99";
			when x"ef" => o_byte <= x"61";
			when x"f0" => o_byte <= x"17";
			when x"f1" => o_byte <= x"2b";
			when x"f2" => o_byte <= x"04";
			when x"f3" => o_byte <= x"7e";
			when x"f4" => o_byte <= x"ba";
			when x"f5" => o_byte <= x"77";
			when x"f6" => o_byte <= x"d6";
			when x"f7" => o_byte <= x"26";
			when x"f8" => o_byte <= x"e1";
			when x"f9" => o_byte <= x"69";
			when x"fa" => o_byte <= x"14";
			when x"fb" => o_byte <= x"63";
			when x"fc" => o_byte <= x"55";
			when x"fd" => o_byte <= x"21";
			when x"fe" => o_byte <= x"0c";
			when x"ff" => o_byte <= x"7d";
			when others => null;
		end case;
	end process;

end architecture behavioral;